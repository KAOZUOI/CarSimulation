// module divider_1ms(input clk, input rst, output reg divided_clk);


module divider_1ms_sim();
    wire clk_s;
    wire rst_s;
    reg divided_clk_s;
    
endmodule